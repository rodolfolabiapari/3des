library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity q_rom is
	port(
		clk 	: IN std_logic;
		address 	: IN std_logic_vector(7 DOWNTO 0);
      data_out : OUT std_logic_vector(3 DOWNTO 0)
	);
end q_rom;

architecture q_rom_behav of q_rom is
type memory is array (integer range 0 to 255) of std_logic_vector (3 downto 0);
  constant mem_Rom : memory := (
	--  q0 t0 0-15
	-- 0X  XX XXXX
	-- 0x8, 0x1, 0x7, 0xd, 0x6, 0xf, 0x3, 0x2, 0x0, 0xb, 0x5, 0x9, 0xe, 0xc, 0xa, 0x4, //00-15
	-- 00000000 a 00001111
			0 => "1000",
			1 => "0001",
			2 => "0111",
			3 => "1101",
			4 => "0110",
			5 => "1111",
			6 => "0011",
			7 => "0010",
			8 => "0000",
			9 => "1011",
			10 => "0101",
			11 => "1001",
			12 => "1110",
			13 => "1100",
			14 => "1010",
			15 => "0100",		
	--  q0 t1 0-15
	-- 0X  XX XXXX
	-- 0xe, 0xc, 0xb, 0x8, 0x1, 0x2, 0x3, 0x5, 0xf, 0x4, 0xa, 0x6, 0x7, 0x0, 0x9, 0xd, //16-31
	-- 00010000 a 00011111
			16 => "1110",
			17 => "1100",
			18 => "1011",
			19 => "1000",
			20 => "0001",
			21 => "0010",
			22 => "0011",
			23 => "0101",
			24 => "1111",
			25 => "0100",
			26 => "1010",
			27 => "0110",
			28 => "0111",
			29 => "0000",
			30 => "1001",
			31 => "1101",		
	--  q0 t2 0-15
	-- 0X  XX XXXX
	-- 0xb, 0xa, 0x5, 0xe, 0x6, 0xd, 0x9, 0x0, 0xc, 0x8, 0xf, 0x3, 0x2, 0x4, 0x7, 0x1, //32-47
	-- 00100000 a 00101111
			32 => "1011",
			33 => "1010",
			34 => "0101",
			35 => "1110",
			36 => "0110",
			37 => "1101",
			38 => "1001",
			39 => "0000",
			40 => "1100",
			41 => "1000",
			42 => "1111",
			43 => "0011",
			44 => "0010",
			45 => "0100",
			46 => "0111",
			47 => "0001",			
	--  q0 t3 0-15
	-- 0X  XX XXXX
	-- 0xd, 0x7, 0xf, 0x4, 0x1, 0x2, 0x6, 0xe, 0x9, 0xb, 0x3, 0x0, 0x8, 0x5, 0xc, 0xa; //48-63
	-- 00110000 a 00111111
			48 => "1101",
			49 => "0111",
			50 => "1111",
			51 => "0100",
			52 => "0001",
			53 => "0010",
			54 => "0110",
			55 => "1110",
			56 => "1001",
			57 => "1011",
			58 => "0011",
			59 => "0000",
			60 => "1000",
			61 => "0101",
			62 => "1100",
			63 => "1010",				
	--  q1 t0 0-15
	-- 0X  XX XXXX
	-- 0x2, 0x8, 0xb, 0xd, 0xf, 0x7, 0x6, 0xe, 0x3, 0x1, 0x9, 0x4, 0x0, 0xa, 0xc, 0x5, //00-15
	-- 01000000 a 01001111
			64 => "0010",
			65 => "1000",
			66 => "1011",
			67 => "1101",
			68 => "1111",
			69 => "0111",
			70 => "0110",
			71 => "1110",
			72 => "0011",
			73 => "0001",
			74 => "1001",
			75 => "0100",
			76 => "0000",
			77 => "1010",
			78 => "1100",
			79 => "0101",	
	--  q1 t1 0-15
	-- 0X  XX XXXX
	-- 0x1, 0xe, 0x2, 0xb, 0x4, 0xc, 0x3, 0x7, 0x6, 0xd, 0xa, 0x5, 0xf, 0x9, 0x0, 0x8, //16-31
	-- 01010000 a 01011111
			80 => "0001",
			81 => "1110",
			82 => "0010",
			83 => "1011",
			84 => "0100",
			85 => "1100",
			86 => "0011",
			87 => "0111",
			88 => "0110",
			89 => "1101",
			90 => "1010",
			91 => "0101",
			92 => "1111",
			93 => "1001",
			94 => "0000",
			95 => "1000",	
	--  q1 t2 0-15
	-- 0X  XX XXXX
	-- 0x4, 0xc, 0x7, 0x5, 0x1, 0x6, 0x9, 0xa, 0x0, 0xe, 0xd, 0x8, 0x2, 0xb, 0x3, 0xf, //32-47
	-- 01100000 a 01101111
			96 => "0100",
			97 => "1100",
			98 => "0111",
			99 => "0101",
			100 => "0001",
			101 => "0110",
			102 => "1001",
			103 => "1010",
			104 => "0000",
			105 => "1110",
			106 => "1101",
			107 => "1000",
			108 => "0010",
			109 => "1011",
			110 => "0011",
			111 => "1111",		
	--  q1 t3 0-15
	-- 0X  XX XXXX
	-- 0xb, 0x9, 0x5, 0x1, 0xc, 0x3, 0xd, 0xe, 0x6, 0x4, 0x7, 0xf, 0x2, 0x0, 0x8, 0xa //48-63
	-- 01110000 a 01111111
			112 => "1011",
			113 => "1001",
			114 => "0101",
			115 => "0001",
			116 => "1100",
			117 => "0011",
			118 => "1101",
			119 => "1110",
			120 => "0110",
			121 => "0100",
			122 => "0111",
			123 => "1111",
			124 => "0010",
			125 => "0000",
			126 => "1000",
			127 => "1010",
	-- 10000000 até 11111111
			others => "0000"
		);
begin
	process(clk)
	begin
		if (clk'event and clk='1') then
			data_out <= mem_Rom(to_integer(unsigned(address)));
		end if;
	end process;
end q_rom_behav;